-- Copyright (C) 1991-2010 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 9.1 Build 350 03/24/2010 Service Pack 2 SJ Full Version"
-- CREATED		"Tue Jun 11 20:17:13 2024"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY dy_time IS 
	PORT
	(
		clk100 :  IN  STD_LOGIC;
		clk10 :  IN  STD_LOGIC;
		clk1 :  IN  STD_LOGIC;
		sel1 :  IN  STD_LOGIC;
		sel2 :  IN  STD_LOGIC;
		sel3 :  IN  STD_LOGIC;
		sel4 :  IN  STD_LOGIC;
		clk1000 :  IN  STD_LOGIC;
		start :  IN  STD_LOGIC;
		sc :  IN  STD_LOGIC;
		clk0_5 :  IN  STD_LOGIC;
		output_A :  OUT  STD_LOGIC;
		output_B :  OUT  STD_LOGIC;
		output_C :  OUT  STD_LOGIC;
		output_D :  OUT  STD_LOGIC;
		output_E :  OUT  STD_LOGIC;
		output_F :  OUT  STD_LOGIC;
		output_G :  OUT  STD_LOGIC;
		end_flag :  OUT  STD_LOGIC;
		fail_flag :  OUT  STD_LOGIC;
		zz :  OUT  STD_LOGIC;
		success :  OUT  STD_LOGIC
	);
END dy_time;

ARCHITECTURE bdf_type OF dy_time IS 

ATTRIBUTE black_box : BOOLEAN;
ATTRIBUTE noopt : BOOLEAN;

COMPONENT \74160_1\
	PORT(CLK : IN STD_LOGIC;
		 ENT : IN STD_LOGIC;
		 LDN : IN STD_LOGIC;
		 ENP : IN STD_LOGIC;
		 QD : OUT STD_LOGIC;
		 QA : OUT STD_LOGIC;
		 QB : OUT STD_LOGIC;
		 QC : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74160_1\: COMPONENT IS true;
ATTRIBUTE noopt OF \74160_1\: COMPONENT IS true;

COMPONENT \74160_2\
	PORT(CLK : IN STD_LOGIC;
		 ENT : IN STD_LOGIC;
		 LDN : IN STD_LOGIC;
		 ENP : IN STD_LOGIC;
		 CLRN : IN STD_LOGIC;
		 QD : OUT STD_LOGIC;
		 QA : OUT STD_LOGIC;
		 QB : OUT STD_LOGIC;
		 QC : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74160_2\: COMPONENT IS true;
ATTRIBUTE noopt OF \74160_2\: COMPONENT IS true;

COMPONENT \74160_6\
	PORT(CLK : IN STD_LOGIC;
		 ENT : IN STD_LOGIC;
		 LDN : IN STD_LOGIC;
		 ENP : IN STD_LOGIC;
		 CLRN : IN STD_LOGIC;
		 QD : OUT STD_LOGIC;
		 QA : OUT STD_LOGIC;
		 QB : OUT STD_LOGIC;
		 QC : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74160_6\: COMPONENT IS true;
ATTRIBUTE noopt OF \74160_6\: COMPONENT IS true;

COMPONENT \74160_7\
	PORT(CLK : IN STD_LOGIC;
		 ENT : IN STD_LOGIC;
		 LDN : IN STD_LOGIC;
		 ENP : IN STD_LOGIC;
		 CLRN : IN STD_LOGIC;
		 QD : OUT STD_LOGIC;
		 QA : OUT STD_LOGIC;
		 QB : OUT STD_LOGIC;
		 QC : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74160_7\: COMPONENT IS true;
ATTRIBUTE noopt OF \74160_7\: COMPONENT IS true;

COMPONENT \74161_0\
	PORT(CLRN : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 ENP : IN STD_LOGIC;
		 LDN : IN STD_LOGIC;
		 A : IN STD_LOGIC;
		 D : IN STD_LOGIC;
		 ENT : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 QD : OUT STD_LOGIC;
		 QC : OUT STD_LOGIC;
		 QB : OUT STD_LOGIC;
		 QA : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74161_0\: COMPONENT IS true;
ATTRIBUTE noopt OF \74161_0\: COMPONENT IS true;

COMPONENT \74244_3\
	PORT(1A2 : IN STD_LOGIC;
		 1A4 : IN STD_LOGIC;
		 1A1 : IN STD_LOGIC;
		 1A3 : IN STD_LOGIC;
		 1GN : IN STD_LOGIC;
		 2A3 : IN STD_LOGIC;
		 2GN : IN STD_LOGIC;
		 2A1 : IN STD_LOGIC;
		 2A4 : IN STD_LOGIC;
		 2A2 : IN STD_LOGIC;
		 1Y2 : OUT STD_LOGIC;
		 1Y4 : OUT STD_LOGIC;
		 2Y1 : OUT STD_LOGIC;
		 1Y1 : OUT STD_LOGIC;
		 2Y3 : OUT STD_LOGIC;
		 2Y4 : OUT STD_LOGIC;
		 1Y3 : OUT STD_LOGIC;
		 2Y2 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74244_3\: COMPONENT IS true;
ATTRIBUTE noopt OF \74244_3\: COMPONENT IS true;

COMPONENT \74244_4\
	PORT(1A2 : IN STD_LOGIC;
		 1A4 : IN STD_LOGIC;
		 1A1 : IN STD_LOGIC;
		 1A3 : IN STD_LOGIC;
		 1GN : IN STD_LOGIC;
		 2A3 : IN STD_LOGIC;
		 2GN : IN STD_LOGIC;
		 2A1 : IN STD_LOGIC;
		 2A4 : IN STD_LOGIC;
		 2A2 : IN STD_LOGIC;
		 1Y2 : OUT STD_LOGIC;
		 1Y4 : OUT STD_LOGIC;
		 2Y1 : OUT STD_LOGIC;
		 1Y1 : OUT STD_LOGIC;
		 2Y3 : OUT STD_LOGIC;
		 2Y4 : OUT STD_LOGIC;
		 1Y3 : OUT STD_LOGIC;
		 2Y2 : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \74244_4\: COMPONENT IS true;
ATTRIBUTE noopt OF \74244_4\: COMPONENT IS true;

COMPONENT \7448_5\
	PORT(A : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 D : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 RBIN : IN STD_LOGIC;
		 BIN : IN STD_LOGIC;
		 LTN : IN STD_LOGIC;
		 OC : OUT STD_LOGIC;
		 OE : OUT STD_LOGIC;
		 OD : OUT STD_LOGIC;
		 OF : OUT STD_LOGIC;
		 OG : OUT STD_LOGIC;
		 OB : OUT STD_LOGIC;
		 OA : OUT STD_LOGIC);
END COMPONENT;
ATTRIBUTE black_box OF \7448_5\: COMPONENT IS true;
ATTRIBUTE noopt OF \7448_5\: COMPONENT IS true;

SIGNAL	SYNTHESIZED_WIRE_71 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_72 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_73 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_74 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_75 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_76 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_77 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_78 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_79 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_80 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_81 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_82 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_83 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_84 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_50 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;
SIGNAL	DFF_inst17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_85 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;


BEGIN 
end_flag <= SYNTHESIZED_WIRE_72;
fail_flag <= SYNTHESIZED_WIRE_51;
zz <= SYNTHESIZED_WIRE_74;
SYNTHESIZED_WIRE_71 <= '1';
SYNTHESIZED_WIRE_6 <= '0';
SYNTHESIZED_WIRE_73 <= '1';
SYNTHESIZED_WIRE_84 <= '1';
SYNTHESIZED_WIRE_85 <= '1';



b2v_inst : 74161_0
PORT MAP(CLRN => start,
		 CLK => clk0_5,
		 ENP => SYNTHESIZED_WIRE_71,
		 LDN => SYNTHESIZED_WIRE_72,
		 A => SYNTHESIZED_WIRE_71,
		 D => SYNTHESIZED_WIRE_71,
		 ENT => SYNTHESIZED_WIRE_71,
		 B => SYNTHESIZED_WIRE_71,
		 C => SYNTHESIZED_WIRE_6,
		 QD => SYNTHESIZED_WIRE_58,
		 QC => SYNTHESIZED_WIRE_61,
		 QB => SYNTHESIZED_WIRE_59,
		 QA => SYNTHESIZED_WIRE_57);



b2v_inst10 : 74160_1
PORT MAP(CLK => clk1000,
		 ENT => SYNTHESIZED_WIRE_72,
		 LDN => SYNTHESIZED_WIRE_73,
		 ENP => sc,
		 QD => SYNTHESIZED_WIRE_78,
		 QA => SYNTHESIZED_WIRE_25,
		 QB => SYNTHESIZED_WIRE_23,
		 QC => SYNTHESIZED_WIRE_26);


b2v_inst11 : 74160_2
PORT MAP(CLK => SYNTHESIZED_WIRE_9,
		 ENT => SYNTHESIZED_WIRE_73,
		 LDN => SYNTHESIZED_WIRE_73,
		 ENP => SYNTHESIZED_WIRE_73,
		 CLRN => SYNTHESIZED_WIRE_74,
		 QD => SYNTHESIZED_WIRE_79,
		 QA => SYNTHESIZED_WIRE_28,
		 QB => SYNTHESIZED_WIRE_30,
		 QC => SYNTHESIZED_WIRE_27);


b2v_inst12 : 74244_3
PORT MAP(1A2 => SYNTHESIZED_WIRE_13,
		 1A4 => SYNTHESIZED_WIRE_75,
		 1A1 => SYNTHESIZED_WIRE_15,
		 1A3 => SYNTHESIZED_WIRE_16,
		 1GN => sel3,
		 2A3 => SYNTHESIZED_WIRE_17,
		 2GN => sel4,
		 2A1 => SYNTHESIZED_WIRE_76,
		 2A4 => SYNTHESIZED_WIRE_19,
		 2A2 => SYNTHESIZED_WIRE_77,
		 1Y2 => SYNTHESIZED_WIRE_83,
		 1Y4 => SYNTHESIZED_WIRE_82,
		 2Y1 => SYNTHESIZED_WIRE_80,
		 1Y1 => SYNTHESIZED_WIRE_80,
		 2Y3 => SYNTHESIZED_WIRE_81,
		 2Y4 => SYNTHESIZED_WIRE_82,
		 1Y3 => SYNTHESIZED_WIRE_81,
		 2Y2 => SYNTHESIZED_WIRE_83);


SYNTHESIZED_WIRE_51 <= SYNTHESIZED_WIRE_77 OR SYNTHESIZED_WIRE_76;


b2v_inst14 : 74244_4
PORT MAP(1A2 => SYNTHESIZED_WIRE_23,
		 1A4 => SYNTHESIZED_WIRE_78,
		 1A1 => SYNTHESIZED_WIRE_25,
		 1A3 => SYNTHESIZED_WIRE_26,
		 1GN => sel1,
		 2A3 => SYNTHESIZED_WIRE_27,
		 2GN => sel2,
		 2A1 => SYNTHESIZED_WIRE_28,
		 2A4 => SYNTHESIZED_WIRE_79,
		 2A2 => SYNTHESIZED_WIRE_30,
		 1Y2 => SYNTHESIZED_WIRE_83,
		 1Y4 => SYNTHESIZED_WIRE_82,
		 2Y1 => SYNTHESIZED_WIRE_80,
		 1Y1 => SYNTHESIZED_WIRE_80,
		 2Y3 => SYNTHESIZED_WIRE_81,
		 2Y4 => SYNTHESIZED_WIRE_82,
		 1Y3 => SYNTHESIZED_WIRE_81,
		 2Y2 => SYNTHESIZED_WIRE_83);


b2v_inst15 : 7448_5
PORT MAP(A => SYNTHESIZED_WIRE_80,
		 C => SYNTHESIZED_WIRE_81,
		 D => SYNTHESIZED_WIRE_82,
		 B => SYNTHESIZED_WIRE_83,
		 RBIN => SYNTHESIZED_WIRE_84,
		 BIN => SYNTHESIZED_WIRE_84,
		 LTN => SYNTHESIZED_WIRE_84,
		 OC => output_C,
		 OE => output_E,
		 OD => output_D,
		 OF => output_F,
		 OG => output_G,
		 OB => output_B,
		 OA => output_A);



PROCESS(SYNTHESIZED_WIRE_50,SYNTHESIZED_WIRE_74)
BEGIN
IF (SYNTHESIZED_WIRE_74 = '0') THEN
	DFF_inst17 <= '1';
ELSIF (RISING_EDGE(SYNTHESIZED_WIRE_50)) THEN
	DFF_inst17 <= SYNTHESIZED_WIRE_51;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_9 <= NOT(SYNTHESIZED_WIRE_78);



SYNTHESIZED_WIRE_63 <= NOT(SYNTHESIZED_WIRE_79);




SYNTHESIZED_WIRE_67 <= NOT(SYNTHESIZED_WIRE_75);



success <= NOT(DFF_inst17);



PROCESS(clk0_5,start,SYNTHESIZED_WIRE_85)
BEGIN
IF (start = '0') THEN
	SYNTHESIZED_WIRE_74 <= '0';
ELSIF (SYNTHESIZED_WIRE_85 = '0') THEN
	SYNTHESIZED_WIRE_74 <= '1';
ELSIF (RISING_EDGE(clk0_5)) THEN
	SYNTHESIZED_WIRE_74 <= SYNTHESIZED_WIRE_85;
END IF;
END PROCESS;



SYNTHESIZED_WIRE_72 <= NOT(SYNTHESIZED_WIRE_57 AND SYNTHESIZED_WIRE_58 AND SYNTHESIZED_WIRE_59 AND SYNTHESIZED_WIRE_60);


SYNTHESIZED_WIRE_60 <= NOT(SYNTHESIZED_WIRE_61);



SYNTHESIZED_WIRE_50 <= NOT(SYNTHESIZED_WIRE_72);



b2v_inst7 : 74160_6
PORT MAP(CLK => SYNTHESIZED_WIRE_63,
		 ENT => SYNTHESIZED_WIRE_73,
		 LDN => SYNTHESIZED_WIRE_73,
		 ENP => SYNTHESIZED_WIRE_73,
		 CLRN => SYNTHESIZED_WIRE_74,
		 QD => SYNTHESIZED_WIRE_75,
		 QA => SYNTHESIZED_WIRE_15,
		 QB => SYNTHESIZED_WIRE_13,
		 QC => SYNTHESIZED_WIRE_16);


b2v_inst8 : 74160_7
PORT MAP(CLK => SYNTHESIZED_WIRE_67,
		 ENT => SYNTHESIZED_WIRE_73,
		 LDN => SYNTHESIZED_WIRE_73,
		 ENP => SYNTHESIZED_WIRE_73,
		 CLRN => SYNTHESIZED_WIRE_74,
		 QD => SYNTHESIZED_WIRE_19,
		 QA => SYNTHESIZED_WIRE_76,
		 QB => SYNTHESIZED_WIRE_77,
		 QC => SYNTHESIZED_WIRE_17);



END bdf_type;